module notgate(input x, output z);


not not1(z,x);
endmodule

