module orgate(input x,input y, output z);


or or1(z,x,y);
endmodule