module andgate(input x,input y, output z);


and and1(z,x,y);
endmodule



