module nandgate(input x,input y, output z);


nand nand1(z,x,y);
endmodule

