module xorgate(input x,input y, output z);


xor xor1(z,x,y);
endmodule